module FSM(IR_15_12, pos, 